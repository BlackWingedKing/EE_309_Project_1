library ieee;

use ieee.std_logic_1164.all;


entity nand16 is

	port(xin,yin: in std_logic_vector(15 downto 0);
		  zout: out std_logic_vector(15 downto 0));

end entity;

architecture arith of nand16 is

begin
	zout(0) <= xin(0) nand yin(0);
	zout(1) <= xin(1) nand yin(1);
	zout(2) <= xin(2) nand yin(2);
	zout(3) <= xin(3) nand yin(3);
	zout(4) <= xin(4) nand yin(4);
	zout(5) <= xin(5) nand yin(5);
	zout(6) <= xin(6) nand yin(6);
	zout(7) <= xin(7) nand yin(7);
	zout(8) <= xin(8) nand yin(8);
	zout(9) <= xin(9) nand yin(9);
	zout(10) <= xin(10) nand yin(10);
	zout(11) <= xin(11) nand yin(11);
	zout(12) <= xin(12) nand yin(12);
	zout(13) <= xin(13) nand yin(13);
	zout(14) <= xin(14) nand yin(14);
	zout(15) <= xin(15) nand yin(15);
end arith;
